module logic2(A, B, Y);
  input A, B;
  output Y;
  or(Y, A, B);
endmodule
