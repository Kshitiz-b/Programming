module logic1(A, B, Y);
  input A, B;
  output Y;
  and(Y, A, B);
endmodule
